architecture pam_map_testbench of TLM_tb is



end architecture pam_map_testbench;