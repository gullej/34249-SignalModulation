-- megafunction wizard: %FIFO%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: dcfifo 

-- ============================================================
-- File Name: clk_sync.vhd
-- Megafunction Name(s):
-- 			dcfifo
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2020  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY clk_sync IS
	GENERIC (
		DATA_WIDTH  : INTEGER);
	PORT
	(
		clk_rd      :  IN  STD_LOGIC;
		clk_wr      :  IN  STD_LOGIC;
		--
		rx_dat      :  IN  STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
		rx_rd       :  IN  STD_LOGIC;
		rx_wr       :  IN  STD_LOGIC;
		--
		tx_dat	    :  OUT STD_LOGIC_VECTOR(8 * DATA_WIDTH - 1 DOWNTO 0);
		tx_empty    :  OUT STD_LOGIC;
		tx_full     :  OUT STD_LOGIC 
	);
END clk_sync;

ARCHITECTURE SYN OF clk_sync IS

	SIGNAL sub_wire0  :  STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
	SIGNAL sub_wire1  :  STD_LOGIC ;
	SIGNAL sub_wire2  :  STD_LOGIC ;

	CONSTANT zeros : STD_LOGIC_VECTOR(7 * DATA_WIDTH - 1 DOWNTO 0) := (others => '0');

	COMPONENT dcfifo
	GENERIC (
		intended_device_family  :  STRING;
		lpm_numwords		    :  NATURAL;
		lpm_showahead		    :  STRING;
		lpm_type		        :  STRING;
		lpm_width		        :  NATURAL;
		lpm_widthu		        :  NATURAL;
		overflow_checking	    :  STRING;
		rdsync_delaypipe	    :  NATURAL;
		underflow_checking	    :  STRING;
		use_eab		            :  STRING;
		wrsync_delaypipe	    :  NATURAL
	);
	PORT (
			data	 :  IN  STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0);
			rdclk	 :  IN  STD_LOGIC ;
			rdreq	 :  IN  STD_LOGIC ;
			wrclk	 :  IN  STD_LOGIC ;
			wrreq	 :  IN  STD_LOGIC ;
			q	     :  OUT STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0);
			rdempty	 :  OUT STD_LOGIC ;
			wrfull	 :  OUT STD_LOGIC 
	); 
	END COMPONENT;

BEGIN
	tx_dat    <= sub_wire0(DATA_WIDTH - 1 DOWNTO 0) & zeros;
	tx_empty  <= sub_wire1;
	tx_full   <= sub_wire2;

	dcfifo_component : dcfifo
	GENERIC MAP (
		intended_device_family => "Cyclone V",
		lpm_numwords           => 32,
		lpm_showahead          => "OFF",
		lpm_type               => "dcfifo",
		lpm_width              => DATA_WIDTH,
		lpm_widthu             => 5,
		overflow_checking      => "ON",
		rdsync_delaypipe       => 5,
		underflow_checking     => "ON",
		use_eab                => "ON",
		wrsync_delaypipe       => 5
	)
	PORT MAP (
		data    => rx_dat,
		rdclk   => clk_rd,
		rdreq   => rx_rd,
		wrclk   => clk_wr,
		wrreq   => rx_wr,
		q       => sub_wire0,
		rdempty => sub_wire1,
		wrfull  => sub_wire2
	);

END SYN;