LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY tranceiver_top IS
    GENERIC (
        DATA_WIDTH : INTEGER);
    PORT (

    );
END tranceiver_top;

ARCHITECTURE tranceiver_top_arc OF tranceiver_top IS
BEGIN

END tranceiver_top_arc;